parameter BIT_WIDTH = 16;